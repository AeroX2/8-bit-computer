--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : computer_fpga                                                ==
--== Component : LogisimToplevelShell                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY LogisimToplevelShell IS
   PORT ( FPGA_INPUT_PIN_0          : IN  std_logic;
          FPGA_INPUT_PIN_1          : IN  std_logic;
          FPGA_OUTPUT_PIN_0         : OUT std_logic;
          FPGA_OUTPUT_PIN_1         : OUT std_logic;
          FPGA_OUTPUT_PIN_2         : OUT std_logic;
          FPGA_OUTPUT_PIN_3         : OUT std_logic;
          FPGA_OUTPUT_PIN_4         : OUT std_logic;
          FPGA_OUTPUT_PIN_5         : OUT std_logic;
          FPGA_OUTPUT_PIN_6         : OUT std_logic;
          FPGA_OUTPUT_PIN_7         : OUT std_logic);
END LogisimToplevelShell;

