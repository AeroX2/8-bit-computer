--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : computer_fpga                                                ==
--== Component : ROM_cu_rom                                                   ==
--==                                                                          ==
--==============================================================================

ARCHITECTURE PlatformIndependent OF ROM_cu_rom IS 

   -----------------------------------------------------------------------------
   -- Here all used signals are defined                                       --
   -----------------------------------------------------------------------------

BEGIN
   MakeRom : PROCESS( Address )
      BEGIN
         CASE (Address) IS
            WHEN "00110000" => Data <= "10000000";
            WHEN "00110001" => Data <= "10000000";
            WHEN "00110010" => Data <= "10000000";
            WHEN "00110011" => Data <= "10000000";
            WHEN "00110100" => Data <= "10000000";
            WHEN "00110101" => Data <= "10000000";
            WHEN "00110110" => Data <= "10000000";
            WHEN "00110111" => Data <= "10000000";
            WHEN "00111000" => Data <= "10000000";
            WHEN "00111001" => Data <= "10000000";
            WHEN "00111010" => Data <= "10000000";
            WHEN "01000000" => Data <= "10000000";
            WHEN "01000001" => Data <= "10000000";
            WHEN "01000010" => Data <= "10000000";
            WHEN "01000011" => Data <= "10000000";
            WHEN "01000100" => Data <= "10000000";
            WHEN "01000101" => Data <= "10000000";
            WHEN "01000110" => Data <= "10000000";
            WHEN "01000111" => Data <= "10000000";
            WHEN "01001000" => Data <= "10000000";
            WHEN "01001001" => Data <= "10000000";
            WHEN "01001010" => Data <= "10000000";
            WHEN "10000000" => Data <= "00100011";
            WHEN "10000001" => Data <= "00100011";
            WHEN "10000010" => Data <= "00100011";
            WHEN "10000011" => Data <= "00110011";
            WHEN "10000100" => Data <= "00110011";
            WHEN "10000101" => Data <= "00110011";
            WHEN "10000110" => Data <= "01000011";
            WHEN "10000111" => Data <= "01000011";
            WHEN "10001000" => Data <= "01000011";
            WHEN "10001001" => Data <= "01010011";
            WHEN "10001010" => Data <= "01010011";
            WHEN "10001011" => Data <= "01010011";
            WHEN "10010011" => Data <= "00100011";
            WHEN "10010100" => Data <= "00110011";
            WHEN "10010101" => Data <= "01000011";
            WHEN "10010110" => Data <= "01010011";
            WHEN "10010111" => Data <= "01010011";
            WHEN "10011000" => Data <= "01010011";
            WHEN OTHERS => Data <= (OTHERS => '0');
         END CASE;
      END PROCESS MakeRom;
END PlatformIndependent;
