--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : computer_fpga                                                ==
--== Component : main                                                         ==
--==                                                                          ==
--==============================================================================


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY main IS
   PORT ( LOGISIM_INPUT_BUBBLES     : IN  std_logic_vector( 0 DOWNTO 0 );
          clk                       : IN  std_logic;
          input_pins                : IN  std_logic_vector( 7 DOWNTO 0 );
          output_pins               : OUT std_logic_vector( 7 DOWNTO 0 ));
END main;

