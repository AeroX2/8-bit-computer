--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : computer_fpga                                                ==
--== Component : ROM_alu_rom                                                  ==
--==                                                                          ==
--==============================================================================

ARCHITECTURE PlatformIndependent OF ROM_alu_rom IS 

   -----------------------------------------------------------------------------
   -- Here all used signals are defined                                       --
   -----------------------------------------------------------------------------

BEGIN
   MakeRom : PROCESS( Address )
      BEGIN
         CASE (Address) IS
            WHEN "00010000" => Data <= "000000100";
            WHEN "00010001" => Data <= "000000100";
            WHEN "00010010" => Data <= "000000001";
            WHEN "00010011" => Data <= "000000001";
            WHEN "00010100" => Data <= "000000001";
            WHEN "00010101" => Data <= "000000001";
            WHEN "00010110" => Data <= "000000101";
            WHEN "00010111" => Data <= "000000101";
            WHEN "00011000" => Data <= "000000101";
            WHEN "00011001" => Data <= "000000101";
            WHEN "00011010" => Data <= "000000101";
            WHEN "00011011" => Data <= "000000101";
            WHEN "00011100" => Data <= "000000101";
            WHEN "00011101" => Data <= "000000101";
            WHEN "00011110" => Data <= "000000101";
            WHEN "00011111" => Data <= "000000101";
            WHEN "00100000" => Data <= "100000100";
            WHEN "00100001" => Data <= "100010010";
            WHEN "00100010" => Data <= "100010010";
            WHEN "00100011" => Data <= "100000001";
            WHEN "00100100" => Data <= "100011000";
            WHEN "00100101" => Data <= "100000000";
            WHEN "00100110" => Data <= "100000001";
            WHEN "00100111" => Data <= "100011000";
            WHEN "00101000" => Data <= "100000000";
            WHEN "01010000" => Data <= "100000101";
            WHEN "01010001" => Data <= "100011111";
            WHEN "01010010" => Data <= "100000111";
            WHEN "01010011" => Data <= "100000100";
            WHEN "01010100" => Data <= "100000001";
            WHEN "01010101" => Data <= "100010100";
            WHEN "01010110" => Data <= "100010001";
            WHEN "01010111" => Data <= "100011100";
            WHEN "01011000" => Data <= "100010011";
            WHEN "01011001" => Data <= "100011110";
            WHEN "01011010" => Data <= "100011011";
            WHEN "01011011" => Data <= "100001100";
            WHEN "01011100" => Data <= "100000011";
            WHEN "01011101" => Data <= "100000000";
            WHEN "01011110" => Data <= "100010010";
            WHEN "01011111" => Data <= "100011000";
            WHEN "01100000" => Data <= "101000000";
            WHEN "01100001" => Data <= "101011010";
            WHEN "01100010" => Data <= "100100000";
            WHEN "01100011" => Data <= "110000000";
            WHEN "01100100" => Data <= "100000101";
            WHEN "01100101" => Data <= "100000101";
            WHEN "01100110" => Data <= "100000101";
            WHEN "01100111" => Data <= "100000101";
            WHEN "01101000" => Data <= "100000101";
            WHEN "01101001" => Data <= "100000101";
            WHEN "01101010" => Data <= "100000101";
            WHEN "01101011" => Data <= "100000101";
            WHEN "01101100" => Data <= "100000101";
            WHEN "01101101" => Data <= "100000101";
            WHEN "01101110" => Data <= "100000101";
            WHEN "01101111" => Data <= "100000101";
            WHEN "10000000" => Data <= "000000100";
            WHEN "10000001" => Data <= "000000100";
            WHEN "10000010" => Data <= "000000100";
            WHEN "10000011" => Data <= "000000001";
            WHEN "10000100" => Data <= "000000001";
            WHEN "10000101" => Data <= "000000001";
            WHEN "10000110" => Data <= "000000001";
            WHEN "10000111" => Data <= "000000001";
            WHEN "10001000" => Data <= "000000001";
            WHEN "10010000" => Data <= "000000100";
            WHEN "10010001" => Data <= "000000001";
            WHEN "10010010" => Data <= "000000001";
            WHEN "10010011" => Data <= "000000100";
            WHEN "10010100" => Data <= "000000001";
            WHEN "10010101" => Data <= "000000001";
            WHEN "10010110" => Data <= "000000100";
            WHEN "10010111" => Data <= "000000001";
            WHEN "10011000" => Data <= "000000001";
            WHEN "10011001" => Data <= "000000100";
            WHEN "10011010" => Data <= "000000001";
            WHEN "10011011" => Data <= "000000001";
            WHEN "10011100" => Data <= "000000100";
            WHEN "10011101" => Data <= "000000001";
            WHEN "10011110" => Data <= "000000001";
            WHEN "10100000" => Data <= "000000101";
            WHEN "10100001" => Data <= "000000101";
            WHEN "10100010" => Data <= "000000101";
            WHEN "10100011" => Data <= "000000101";
            WHEN "10100100" => Data <= "000000101";
            WHEN "10100101" => Data <= "000000101";
            WHEN "10110000" => Data <= "000000100";
            WHEN "10110001" => Data <= "000000001";
            WHEN "10110010" => Data <= "000000001";
            WHEN "11000000" => Data <= "000000100";
            WHEN "11000001" => Data <= "000000001";
            WHEN "11000010" => Data <= "000000001";
            WHEN OTHERS => Data <= (OTHERS => '0');
         END CASE;
      END PROCESS MakeRom;
END PlatformIndependent;
