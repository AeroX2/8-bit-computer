--==============================================================================
--== Logisim goes FPGA automatic generated VHDL code                          ==
--==                                                                          ==
--==                                                                          ==
--== Project   : computer_fpga                                                ==
--== Component : ROM_cu_rom_2                                                 ==
--==                                                                          ==
--==============================================================================

ARCHITECTURE PlatformIndependent OF ROM_cu_rom_2 IS 

   -----------------------------------------------------------------------------
   -- Here all used signals are defined                                       --
   -----------------------------------------------------------------------------

BEGIN
   MakeRom : PROCESS( Address )
      BEGIN
         CASE (Address) IS
            WHEN "00010000" => Data <= "00100101";
            WHEN "00010001" => Data <= "00100110";
            WHEN "00010010" => Data <= "00110100";
            WHEN "00010011" => Data <= "00100110";
            WHEN "00010100" => Data <= "01000100";
            WHEN "00010101" => Data <= "01000101";
            WHEN "00100000" => Data <= "00100000";
            WHEN "00100001" => Data <= "00100000";
            WHEN "00100010" => Data <= "01000000";
            WHEN "00100011" => Data <= "00100000";
            WHEN "00100100" => Data <= "00100000";
            WHEN "00100110" => Data <= "01000000";
            WHEN "00100111" => Data <= "01000000";
            WHEN "00110000" => Data <= "11110000";
            WHEN "00110001" => Data <= "11110000";
            WHEN "00110010" => Data <= "11110000";
            WHEN "00110011" => Data <= "11110000";
            WHEN "00110100" => Data <= "11110000";
            WHEN "00110101" => Data <= "11110000";
            WHEN "00110110" => Data <= "11110000";
            WHEN "00110111" => Data <= "11110000";
            WHEN "00111000" => Data <= "11110000";
            WHEN "00111001" => Data <= "11110000";
            WHEN "00111010" => Data <= "11110000";
            WHEN "01000000" => Data <= "11110000";
            WHEN "01000001" => Data <= "11110000";
            WHEN "01000010" => Data <= "11110000";
            WHEN "01000011" => Data <= "11110000";
            WHEN "01000100" => Data <= "11110000";
            WHEN "01000101" => Data <= "11110000";
            WHEN "01000110" => Data <= "11110000";
            WHEN "01000111" => Data <= "11110000";
            WHEN "01001000" => Data <= "11110000";
            WHEN "01001001" => Data <= "11110000";
            WHEN "01001010" => Data <= "11110000";
            WHEN "01010000" => Data <= "00110100";
            WHEN "01010001" => Data <= "00110100";
            WHEN "01010010" => Data <= "00110100";
            WHEN "01010011" => Data <= "00110100";
            WHEN "01010100" => Data <= "00110100";
            WHEN "01010101" => Data <= "00110100";
            WHEN "01010110" => Data <= "00110100";
            WHEN "01010111" => Data <= "00110100";
            WHEN "01011000" => Data <= "00110100";
            WHEN "01011001" => Data <= "00110100";
            WHEN "01011010" => Data <= "00110100";
            WHEN "01011011" => Data <= "00110100";
            WHEN "01011100" => Data <= "00110100";
            WHEN "01011101" => Data <= "00110100";
            WHEN "01011110" => Data <= "00110100";
            WHEN "01011111" => Data <= "00110100";
            WHEN "01100000" => Data <= "00110100";
            WHEN "01100001" => Data <= "00110100";
            WHEN "01100010" => Data <= "00110100";
            WHEN "01100011" => Data <= "00110100";
            WHEN "01100100" => Data <= "00110100";
            WHEN "01100101" => Data <= "00110100";
            WHEN "01100110" => Data <= "00110100";
            WHEN "01100111" => Data <= "00110100";
            WHEN "01101000" => Data <= "00110100";
            WHEN "01101001" => Data <= "00110100";
            WHEN "01101010" => Data <= "00110100";
            WHEN "01101011" => Data <= "00110100";
            WHEN "01101100" => Data <= "00110100";
            WHEN "01101101" => Data <= "00110100";
            WHEN "01101110" => Data <= "00110100";
            WHEN "01101111" => Data <= "00110100";
            WHEN "01110000" => Data <= "11010100";
            WHEN "01110001" => Data <= "11010101";
            WHEN "01110010" => Data <= "11010110";
            WHEN "10000000" => Data <= "01100100";
            WHEN "10000001" => Data <= "01100101";
            WHEN "10000010" => Data <= "01100110";
            WHEN "10000011" => Data <= "01100100";
            WHEN "10000100" => Data <= "01100101";
            WHEN "10000101" => Data <= "01100110";
            WHEN "10000110" => Data <= "01100100";
            WHEN "10000111" => Data <= "01100101";
            WHEN "10001000" => Data <= "01100110";
            WHEN "10001001" => Data <= "01100100";
            WHEN "10001010" => Data <= "01100101";
            WHEN "10001011" => Data <= "01100110";
            WHEN "10010000" => Data <= "00100010";
            WHEN "10010001" => Data <= "00110010";
            WHEN "10010010" => Data <= "01000010";
            WHEN "10010011" => Data <= "00100010";
            WHEN "10010100" => Data <= "00110010";
            WHEN "10010101" => Data <= "01000010";
            WHEN "10010110" => Data <= "00100010";
            WHEN "10010111" => Data <= "00110010";
            WHEN "10011000" => Data <= "01000010";
            WHEN "10011001" => Data <= "00100011";
            WHEN "10011010" => Data <= "00110011";
            WHEN "10011011" => Data <= "01000011";
            WHEN "10100000" => Data <= "00010100";
            WHEN "10100001" => Data <= "00010101";
            WHEN "10100010" => Data <= "00010110";
            WHEN "10110000" => Data <= "00100001";
            WHEN "10110001" => Data <= "00110001";
            WHEN "10110010" => Data <= "01000001";
            WHEN "11110000" => Data <= "00001111";
            WHEN OTHERS => Data <= (OTHERS => '0');
         END CASE;
      END PROCESS MakeRom;
END PlatformIndependent;
